module ShiftRows_tb();
 reg [127 : 0 ] in;
 wire  [127 : 0 ] out ;

initial begin
in = 128'h_adcb0f257e9c63e0bc557e951c15ef01;
# 50;
in = 128'h_884a33781fdb75c2d380349e19f876fb;  
end



ShiftRows ShiftRows_dut(
    .in(in),
    .out(out)
);

always @ (in) begin
    $display("in = %h", in);
    $display("out = %h", out);

end

endmodule