module SubByte(stateIn,stateOut);

	input[127:0]stateIn;
	output [127:0]stateOut;
	assign stateOut = stateIn;

endmodule