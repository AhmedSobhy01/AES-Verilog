module SBox(in, out);
    input [7:0] in;
    output [7:0] out;

    reg [7:0] tmp;
    assign out = tmp;

    always @(in) begin
        case (in)
            8'h00: tmp = 8'h63;
            8'h01: tmp = 8'h7c;
            8'h02: tmp = 8'h77;
            8'h03: tmp = 8'h7b;
            8'h04: tmp = 8'hf2;
            8'h05: tmp = 8'h6b;
            8'h06: tmp = 8'h6f;
            8'h07: tmp = 8'hc5;
            8'h08: tmp = 8'h30;
            8'h09: tmp = 8'h01;
            8'h0a: tmp = 8'h67;
            8'h0b: tmp = 8'h2b;
            8'h0c: tmp = 8'hfe;
            8'h0d: tmp = 8'hd7;
            8'h0e: tmp = 8'hab;
            8'h0f: tmp = 8'h76;
            8'h10: tmp = 8'hca;
            8'h11: tmp = 8'h82;
            8'h12: tmp = 8'hc9;
            8'h13: tmp = 8'h7d;
            8'h14: tmp = 8'hfa;
            8'h15: tmp = 8'h59;
            8'h16: tmp = 8'h47;
            8'h17: tmp = 8'hf0;
            8'h18: tmp = 8'had;
            8'h19: tmp = 8'hd4;
            8'h1a: tmp = 8'ha2;
            8'h1b: tmp = 8'haf;
            8'h1c: tmp = 8'h9c;
            8'h1d: tmp = 8'ha4;
            8'h1e: tmp = 8'h72;
            8'h1f: tmp = 8'hc0;
            8'h20: tmp = 8'hb7;
            8'h21: tmp = 8'hfd;
            8'h22: tmp = 8'h93;
            8'h23: tmp = 8'h26;
            8'h24: tmp = 8'h36;
            8'h25: tmp = 8'h3f;
            8'h26: tmp = 8'hf7;
            8'h27: tmp = 8'hcc;
            8'h28: tmp = 8'h34;
            8'h29: tmp = 8'ha5;
            8'h2a: tmp = 8'he5;
            8'h2b: tmp = 8'hf1;
            8'h2c: tmp = 8'h71;
            8'h2d: tmp = 8'hd8;
            8'h2e: tmp = 8'h31;
            8'h2f: tmp = 8'h15;
            8'h30: tmp = 8'h04;
            8'h31: tmp = 8'hc7;
            8'h32: tmp = 8'h23;
            8'h33: tmp = 8'hc3;
            8'h34: tmp = 8'h18;
            8'h35: tmp = 8'h96;
            8'h36: tmp = 8'h05;
            8'h37: tmp = 8'h9a;
            8'h38: tmp = 8'h07;
            8'h39: tmp = 8'h12;
            8'h3a: tmp = 8'h80;
            8'h3b: tmp = 8'he2;
            8'h3c: tmp = 8'heb;
            8'h3d: tmp = 8'h27;
            8'h3e: tmp = 8'hb2;
            8'h3f: tmp = 8'h75;
            8'h40: tmp = 8'h09;
            8'h41: tmp = 8'h83;
            8'h42: tmp = 8'h2c;
            8'h43: tmp = 8'h1a;
            8'h44: tmp = 8'h1b;
            8'h45: tmp = 8'h6e;
            8'h46: tmp = 8'h5a;
            8'h47: tmp = 8'ha0;
            8'h48: tmp = 8'h52;
            8'h49: tmp = 8'h3b;
            8'h4a: tmp = 8'hd6;
            8'h4b: tmp = 8'hb3;
            8'h4c: tmp = 8'h29;
            8'h4d: tmp = 8'he3;
            8'h4e: tmp = 8'h2f;
            8'h4f: tmp = 8'h84;
            8'h50: tmp = 8'h53;
            8'h51: tmp = 8'hd1;
            8'h52: tmp = 8'h00;
            8'h53: tmp = 8'hed;
            8'h54: tmp = 8'h20;
            8'h55: tmp = 8'hfc;
            8'h56: tmp = 8'hb1;
            8'h57: tmp = 8'h5b;
            8'h58: tmp = 8'h6a;
            8'h59: tmp = 8'hcb;
            8'h5a: tmp = 8'hbe;
            8'h5b: tmp = 8'h39;
            8'h5c: tmp = 8'h4a;
            8'h5d: tmp = 8'h4c;
            8'h5e: tmp = 8'h58;
            8'h5f: tmp = 8'hcf;
            8'h60: tmp = 8'hd0;
            8'h61: tmp = 8'hef;
            8'h62: tmp = 8'haa;
            8'h63: tmp = 8'hfb;
            8'h64: tmp = 8'h43;
            8'h65: tmp = 8'h4d;
            8'h66: tmp = 8'h33;
            8'h67: tmp = 8'h85;
            8'h68: tmp = 8'h45;
            8'h69: tmp = 8'hf9;
            8'h6a: tmp = 8'h02;
            8'h6b: tmp = 8'h7f;
            8'h6c: tmp = 8'h50;
            8'h6d: tmp = 8'h3c;
            8'h6e: tmp = 8'h9f;
            8'h6f: tmp = 8'ha8;
            8'h70: tmp = 8'h51;
            8'h71: tmp = 8'ha3;
            8'h72: tmp = 8'h40;
            8'h73: tmp = 8'h8f;
            8'h74: tmp = 8'h92;
            8'h75: tmp = 8'h9d;
            8'h76: tmp = 8'h38;
            8'h77: tmp = 8'hf5;
            8'h78: tmp = 8'hbc;
            8'h79: tmp = 8'hb6;
            8'h7a: tmp = 8'hda;
            8'h7b: tmp = 8'h21;
            8'h7c: tmp = 8'h10;
            8'h7d: tmp = 8'hff;
            8'h7e: tmp = 8'hf3;
            8'h7f: tmp = 8'hd2;
            8'h80: tmp = 8'hcd;
            8'h81: tmp = 8'h0c;
            8'h82: tmp = 8'h13;
            8'h83: tmp = 8'hec;
            8'h84: tmp = 8'h5f;
            8'h85: tmp = 8'h97;
            8'h86: tmp = 8'h44;
            8'h87: tmp = 8'h17;
            8'h88: tmp = 8'hc4;
            8'h89: tmp = 8'ha7;
            8'h8a: tmp = 8'h7e;
            8'h8b: tmp = 8'h3d;
            8'h8c: tmp = 8'h64;
            8'h8d: tmp = 8'h5d;
            8'h8e: tmp = 8'h19;
            8'h8f: tmp = 8'h73;
            8'h90: tmp = 8'h60;
            8'h91: tmp = 8'h81;
            8'h92: tmp = 8'h4f;
            8'h93: tmp = 8'hdc;
            8'h94: tmp = 8'h22;
            8'h95: tmp = 8'h2a;
            8'h96: tmp = 8'h90;
            8'h97: tmp = 8'h88;
            8'h98: tmp = 8'h46;
            8'h99: tmp = 8'hee;
            8'h9a: tmp = 8'hb8;
            8'h9b: tmp = 8'h14;
            8'h9c: tmp = 8'hde;
            8'h9d: tmp = 8'h5e;
            8'h9e: tmp = 8'h0b;
            8'h9f: tmp = 8'hdb;
            8'ha0: tmp = 8'he0;
            8'ha1: tmp = 8'h32;
            8'ha2: tmp = 8'h3a;
            8'ha3: tmp = 8'h0a;
            8'ha4: tmp = 8'h49;
            8'ha5: tmp = 8'h06;
            8'ha6: tmp = 8'h24;
            8'ha7: tmp = 8'h5c;
            8'ha8: tmp = 8'hc2;
            8'ha9: tmp = 8'hd3;
            8'haa: tmp = 8'hac;
            8'hab: tmp = 8'h62;
            8'hac: tmp = 8'h91;
            8'had: tmp = 8'h95;
            8'hae: tmp = 8'he4;
            8'haf: tmp = 8'h79;
            8'hb0: tmp = 8'he7;
            8'hb1: tmp = 8'hc8;
            8'hb2: tmp = 8'h37;
            8'hb3: tmp = 8'h6d;
            8'hb4: tmp = 8'h8d;
            8'hb5: tmp = 8'hd5;
            8'hb6: tmp = 8'h4e;
            8'hb7: tmp = 8'ha9;
            8'hb8: tmp = 8'h6c;
            8'hb9: tmp = 8'h56;
            8'hba: tmp = 8'hf4;
            8'hbb: tmp = 8'hea;
            8'hbc: tmp = 8'h65;
            8'hbd: tmp = 8'h7a;
            8'hbe: tmp = 8'hae;
            8'hbf: tmp = 8'h08;
            8'hc0: tmp = 8'hba;
            8'hc1: tmp = 8'h78;
            8'hc2: tmp = 8'h25;
            8'hc3: tmp = 8'h2e;
            8'hc4: tmp = 8'h1c;
            8'hc5: tmp = 8'ha6;
            8'hc6: tmp = 8'hb4;
            8'hc7: tmp = 8'hc6;
            8'hc8: tmp = 8'he8;
            8'hc9: tmp = 8'hdd;
            8'hca: tmp = 8'h74;
            8'hcb: tmp = 8'h1f;
            8'hcc: tmp = 8'h4b;
            8'hcd: tmp = 8'hbd;
            8'hce: tmp = 8'h8b;
            8'hcf: tmp = 8'h8a;
            8'hd0: tmp = 8'h70;
            8'hd1: tmp = 8'h3e;
            8'hd2: tmp = 8'hb5;
            8'hd3: tmp = 8'h66;
            8'hd4: tmp = 8'h48;
            8'hd5: tmp = 8'h03;
            8'hd6: tmp = 8'hf6;
            8'hd7: tmp = 8'h0e;
            8'hd8: tmp = 8'h61;
            8'hd9: tmp = 8'h35;
            8'hda: tmp = 8'h57;
            8'hdb: tmp = 8'hb9;
            8'hdc: tmp = 8'h86;
            8'hdd: tmp = 8'hc1;
            8'hde: tmp = 8'h1d;
            8'hdf: tmp = 8'h9e;
            8'he0: tmp = 8'he1;
            8'he1: tmp = 8'hf8;
            8'he2: tmp = 8'h98;
            8'he3: tmp = 8'h11;
            8'he4: tmp = 8'h69;
            8'he5: tmp = 8'hd9;
            8'he6: tmp = 8'h8e;
            8'he7: tmp = 8'h94;
            8'he8: tmp = 8'h9b;
            8'he9: tmp = 8'h1e;
            8'hea: tmp = 8'h87;
            8'heb: tmp = 8'he9;
            8'hec: tmp = 8'hce;
            8'hed: tmp = 8'h55;
            8'hee: tmp = 8'h28;
            8'hef: tmp = 8'hdf;
            8'hf0: tmp = 8'h8c;
            8'hf1: tmp = 8'ha1;
            8'hf2: tmp = 8'h89;
            8'hf3: tmp = 8'h0d;
            8'hf4: tmp = 8'hbf;
            8'hf5: tmp = 8'he6;
            8'hf6: tmp = 8'h42;
            8'hf7: tmp = 8'h68;
            8'hf8: tmp = 8'h41;
            8'hf9: tmp = 8'h99;
            8'hfa: tmp = 8'h2d;
            8'hfb: tmp = 8'h0f;
            8'hfc: tmp = 8'hb0;
            8'hfd: tmp = 8'h54;
            8'hfe: tmp = 8'hbb;
            8'hff: tmp = 8'h16;
        endcase
    end
endmodule