module InvShiftRows_tb();
 reg [127 : 0 ] in;
 wire  [127 : 0 ] out ;

initial begin
in = 128'h_aa5ece06ee6e3c56dde68bac2621bebf;
# 50;
in = 128'h_d1ed44fd1a0f3f2afa4ff27b7c332a69;  
end



InvShiftRows InvShiftRows_dut(
    .in(in),
    .out(out)
);

always @ (in) begin
    $display("in = %h", in);
    $display("out = %h", out);

end

endmodule