module InvSubTable(subByte, oriByte);
	input [7:0] subByte; 
	output reg [7:0] oriByte;

	always @(*) begin  
		case (subByte)
			8'h00: oriByte =8'h52;
			8'h01: oriByte =8'h09;
			8'h02: oriByte =8'h6a;
			8'h03: oriByte =8'hd5;
			8'h04: oriByte =8'h30;
			8'h05: oriByte =8'h36;
			8'h06: oriByte =8'ha5;
			8'h07: oriByte =8'h38;
			8'h08: oriByte =8'hbf;
			8'h09: oriByte =8'h40;
			8'h0a: oriByte =8'ha3;
			8'h0b: oriByte =8'h9e;
			8'h0c: oriByte =8'h81;
			8'h0d: oriByte =8'hf3;
			8'h0e: oriByte =8'hd7;
			8'h0f: oriByte =8'hfb;
			8'h10: oriByte =8'h7c;
			8'h11: oriByte =8'he3;
			8'h12: oriByte =8'h39;
			8'h13: oriByte =8'h82;
			8'h14: oriByte =8'h9b;
			8'h15: oriByte =8'h2f;
			8'h16: oriByte =8'hff;
			8'h17: oriByte =8'h87;
			8'h18: oriByte =8'h34;
			8'h19: oriByte =8'h8e;
			8'h1a: oriByte =8'h43;
			8'h1b: oriByte =8'h44;
			8'h1c: oriByte =8'hc4;
			8'h1d: oriByte =8'hde;
			8'h1e: oriByte =8'he9;
			8'h1f: oriByte =8'hcb;
			8'h20: oriByte =8'h54;
			8'h21: oriByte =8'h7b;
			8'h22: oriByte =8'h94;
			8'h23: oriByte =8'h32;
			8'h24: oriByte =8'ha6;
			8'h25: oriByte =8'hc2;
			8'h26: oriByte =8'h23;
			8'h27: oriByte =8'h3d;
			8'h28: oriByte =8'hee;
			8'h29: oriByte =8'h4c;
			8'h2a: oriByte =8'h95;
			8'h2b: oriByte =8'h0b;
			8'h2c: oriByte =8'h42;
			8'h2d: oriByte =8'hfa;
			8'h2e: oriByte =8'hc3;
			8'h2f: oriByte =8'h4e;
			8'h30: oriByte =8'h08;
			8'h31: oriByte =8'h2e;
			8'h32: oriByte =8'ha1;
			8'h33: oriByte =8'h66;
			8'h34: oriByte =8'h28;
			8'h35: oriByte =8'hd9;
			8'h36: oriByte =8'h24;
			8'h37: oriByte =8'hb2;
			8'h38: oriByte =8'h76;
			8'h39: oriByte =8'h5b;
			8'h3a: oriByte =8'ha2;
			8'h3b: oriByte =8'h49;
			8'h3c: oriByte =8'h6d;
			8'h3d: oriByte =8'h8b;
			8'h3e: oriByte =8'hd1;
			8'h3f: oriByte =8'h25;
			8'h40: oriByte =8'h72;
			8'h41: oriByte =8'hf8;
			8'h42: oriByte =8'hf6;
			8'h43: oriByte =8'h64;
			8'h44: oriByte =8'h86;
			8'h45: oriByte =8'h68;
			8'h46: oriByte =8'h98;
			8'h47: oriByte =8'h16;
			8'h48: oriByte =8'hd4;
			8'h49: oriByte =8'ha4;
			8'h4a: oriByte =8'h5c;
			8'h4b: oriByte =8'hcc;
			8'h4c: oriByte =8'h5d;
			8'h4d: oriByte =8'h65;
			8'h4e: oriByte =8'hb6;
			8'h4f: oriByte =8'h92;
			8'h50: oriByte =8'h6c;
			8'h51: oriByte =8'h70;
			8'h52: oriByte =8'h48;
			8'h53: oriByte =8'h50;
			8'h54: oriByte =8'hfd;
			8'h55: oriByte =8'hed;
			8'h56: oriByte =8'hb9;
			8'h57: oriByte =8'hda;
			8'h58: oriByte =8'h5e;
			8'h59: oriByte =8'h15;
			8'h5a: oriByte =8'h46;
			8'h5b: oriByte =8'h57;
			8'h5c: oriByte =8'ha7;
			8'h5d: oriByte =8'h8d;
			8'h5e: oriByte =8'h9d;
			8'h5f: oriByte =8'h84;
			8'h60: oriByte =8'h90;
			8'h61: oriByte =8'hd8;
			8'h62: oriByte =8'hab;
			8'h63: oriByte =8'h00;
			8'h64: oriByte =8'h8c;
			8'h65: oriByte =8'hbc;
			8'h66: oriByte =8'hd3;
			8'h67: oriByte =8'h0a;
			8'h68: oriByte =8'hf7;
			8'h69: oriByte =8'he4;
			8'h6a: oriByte =8'h58;
			8'h6b: oriByte =8'h05;
			8'h6c: oriByte =8'hb8;
			8'h6d: oriByte =8'hb3;
			8'h6e: oriByte =8'h45;
			8'h6f: oriByte =8'h06;
			8'h70: oriByte =8'hd0;
			8'h71: oriByte =8'h2c;
			8'h72: oriByte =8'h1e;
			8'h73: oriByte =8'h8f;
			8'h74: oriByte =8'hca;
			8'h75: oriByte =8'h3f;
			8'h76: oriByte =8'h0f;
			8'h77: oriByte =8'h02;
			8'h78: oriByte =8'hc1;
			8'h79: oriByte =8'haf;
			8'h7a: oriByte =8'hbd;
			8'h7b: oriByte =8'h03;
			8'h7c: oriByte =8'h01;
			8'h7d: oriByte =8'h13;
			8'h7e: oriByte =8'h8a;
			8'h7f: oriByte =8'h6b;
			8'h80: oriByte =8'h3a;
			8'h81: oriByte =8'h91;
			8'h82: oriByte =8'h11;
			8'h83: oriByte =8'h41;
			8'h84: oriByte =8'h4f;
			8'h85: oriByte =8'h67;
			8'h86: oriByte =8'hdc;
			8'h87: oriByte =8'hea;
			8'h88: oriByte =8'h97;
			8'h89: oriByte =8'hf2;
			8'h8a: oriByte =8'hcf;
			8'h8b: oriByte =8'hce;
			8'h8c: oriByte =8'hf0;
			8'h8d: oriByte =8'hb4;
			8'h8e: oriByte =8'he6;
			8'h8f: oriByte =8'h73;
			8'h90: oriByte =8'h96;
			8'h91: oriByte =8'hac;
			8'h92: oriByte =8'h74;
			8'h93: oriByte =8'h22;
			8'h94: oriByte =8'he7;
			8'h95: oriByte =8'had;
			8'h96: oriByte =8'h35;
			8'h97: oriByte =8'h85;
			8'h98: oriByte =8'he2;
			8'h99: oriByte =8'hf9;
			8'h9a: oriByte =8'h37;
			8'h9b: oriByte =8'he8;
			8'h9c: oriByte =8'h1c;
			8'h9d: oriByte =8'h75;
			8'h9e: oriByte =8'hdf;
			8'h9f: oriByte =8'h6e;
			8'ha0: oriByte =8'h47;
			8'ha1: oriByte =8'hf1;
			8'ha2: oriByte =8'h1a;
			8'ha3: oriByte =8'h71;
			8'ha4: oriByte =8'h1d;
			8'ha5: oriByte =8'h29;
			8'ha6: oriByte =8'hc5;
			8'ha7: oriByte =8'h89;
			8'ha8: oriByte =8'h6f;
			8'ha9: oriByte =8'hb7;
			8'haa: oriByte =8'h62;
			8'hab: oriByte =8'h0e;
			8'hac: oriByte =8'haa;
			8'had: oriByte =8'h18;
			8'hae: oriByte =8'hbe;
			8'haf: oriByte =8'h1b;
			8'hb0: oriByte =8'hfc;
			8'hb1: oriByte =8'h56;
			8'hb2: oriByte =8'h3e;
			8'hb3: oriByte =8'h4b;
			8'hb4: oriByte =8'hc6;
			8'hb5: oriByte =8'hd2;
			8'hb6: oriByte =8'h79;
			8'hb7: oriByte =8'h20;
			8'hb8: oriByte =8'h9a;
			8'hb9: oriByte =8'hdb;
			8'hba: oriByte =8'hc0;
			8'hbb: oriByte =8'hfe;
			8'hbc: oriByte =8'h78;
			8'hbd: oriByte =8'hcd;
			8'hbe: oriByte =8'h5a;
			8'hbf: oriByte =8'hf4;
			8'hc0: oriByte =8'h1f;
			8'hc1: oriByte =8'hdd;
			8'hc2: oriByte =8'ha8;
			8'hc3: oriByte =8'h33;
			8'hc4: oriByte =8'h88;
			8'hc5: oriByte =8'h07;
			8'hc6: oriByte =8'hc7;
			8'hc7: oriByte =8'h31;
			8'hc8: oriByte =8'hb1;
			8'hc9: oriByte =8'h12;
			8'hca: oriByte =8'h10;
			8'hcb: oriByte =8'h59;
			8'hcc: oriByte =8'h27;
			8'hcd: oriByte =8'h80;
			8'hce: oriByte =8'hec;
			8'hcf: oriByte =8'h5f;
			8'hd0: oriByte =8'h60;
			8'hd1: oriByte =8'h51;
			8'hd2: oriByte =8'h7f;
			8'hd3: oriByte =8'ha9;
			8'hd4: oriByte =8'h19;
			8'hd5: oriByte =8'hb5;
			8'hd6: oriByte =8'h4a;
			8'hd7: oriByte =8'h0d;
			8'hd8: oriByte =8'h2d;
			8'hd9: oriByte =8'he5;
			8'hda: oriByte =8'h7a;
			8'hdb: oriByte =8'h9f;
			8'hdc: oriByte =8'h93;
			8'hdd: oriByte =8'hc9;
			8'hde: oriByte =8'h9c;
			8'hdf: oriByte =8'hef;
			8'he0: oriByte =8'ha0;
			8'he1: oriByte =8'he0;
			8'he2: oriByte =8'h3b;
			8'he3: oriByte =8'h4d;
			8'he4: oriByte =8'hae;
			8'he5: oriByte =8'h2a;
			8'he6: oriByte =8'hf5;
			8'he7: oriByte =8'hb0;
			8'he8: oriByte =8'hc8;
			8'he9: oriByte =8'heb;
			8'hea: oriByte =8'hbb;
			8'heb: oriByte =8'h3c;
			8'hec: oriByte =8'h83;
			8'hed: oriByte =8'h53;
			8'hee: oriByte =8'h99;
			8'hef: oriByte =8'h61;
			8'hf0: oriByte =8'h17;
			8'hf1: oriByte =8'h2b;
			8'hf2: oriByte =8'h04;
			8'hf3: oriByte =8'h7e;
			8'hf4: oriByte =8'hba;
			8'hf5: oriByte =8'h77;
			8'hf6: oriByte =8'hd6;
			8'hf7: oriByte =8'h26;
			8'hf8: oriByte =8'he1;
			8'hf9: oriByte =8'h69;
			8'hfa: oriByte =8'h14;
			8'hfb: oriByte =8'h63;
			8'hfc: oriByte =8'h55;
			8'hfd: oriByte =8'h21;
			8'hfe: oriByte =8'h0c;
			8'hff: oriByte =8'h7d;
		endcase
	end
endmodule
